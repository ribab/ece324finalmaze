
module maze_carver
	(
		input clk,
		input start,
		input wire [2:0] x_dimension,
		input wire [2:0] y_dimension,
		output reg [64*64-1:0] maze_data,
		output reg finish
	);
	
//	reg [64-1:0] maze_paths [64-1:0];
	
//	 maze_paths
//  000...0
//  111...0
//  000...0
//  ...
//  000...0

	
	reg [15:0] i;
	reg [15:0] j;

	initial begin
		for (i = 0; i < 64; i = i + 1)
			for (j = 0; j < 64; j = j + 1)
				maze_data [i + 64*j] = 0;
		maze_data = 4095'b101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100;
		
	end
	
endmodule
/*
      maze_paths [0] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [1] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [2] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [3] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [4] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [5] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [6] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [7] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [8] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [9] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [10] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [11] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [12] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [13] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [14] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [15] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [16] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [17] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [18] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [19] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [20] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [21] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [22] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [23] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [24] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [25] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [26] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [27] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [28] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [29] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [30] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [31] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [32] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [33] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [34] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [35] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [36] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [37] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [38] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [39] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [40] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [41] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [42] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [43] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [44] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [45] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [46] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [47] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [48] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [49] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [50] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [51] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [52] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [53] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [54] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [55] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [56] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [57] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [58] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [59] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [60] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [61] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [62] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [63] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [64] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [65] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [66] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [67] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [68] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [69] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [70] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [71] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [72] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [73] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [74] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [75] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [76] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [77] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [78] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [79] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [80] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [81] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [82] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [83] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [84] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [85] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [86] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [87] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [88] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [89] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [90] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [91] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [92] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [93] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [94] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [95] = 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [96] = 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [97] = 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [98] = 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [99] = 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
	end
	
	assign maze_data[99:0]     = maze_paths[0];
	assign maze_data[199:100]  = maze_paths[1];
	assign maze_data[299:200]  = maze_paths[2];
	assign maze_data[399:300]  = maze_paths[3];
	assign maze_data[499:400]  = maze_paths[4];
	assign maze_data[599:500]  = maze_paths[5];
	assign maze_data[699:600]  = maze_paths[6];
	assign maze_data[799:700]  = maze_paths[7];
	assign maze_data[899:800]  = maze_paths[8];
	assign maze_data[999:900]  = maze_paths[9];
	assign maze_data[1099:1000]   = maze_paths[10];
	assign maze_data[1199:1100] = maze_paths[11];
	assign maze_data[1299:1200] = maze_paths[12];
	assign maze_data[1399:1300] = maze_paths[13];
	assign maze_data[1499:1400] = maze_paths[14];
	assign maze_data[1599:1500] = maze_paths[15];
	assign maze_data[1699:1600] = maze_paths[16];
	assign maze_data[1799:1700] = maze_paths[17];
	assign maze_data[1899:1800] = maze_paths[18];
	assign maze_data[1999:1900] = maze_paths[19];
	assign maze_data[2099:2000]   = maze_paths[20];
	assign maze_data[2199:2100] = maze_paths[21];
	assign maze_data[2299:2200] = maze_paths[22];
	assign maze_data[2399:2300] = maze_paths[23];
	assign maze_data[2499:2400] = maze_paths[24];
	assign maze_data[2599:2500] = maze_paths[25];
	assign maze_data[2699:2600] = maze_paths[26];
	assign maze_data[2799:2700] = maze_paths[27];
	assign maze_data[2899:2800] = maze_paths[28];
	assign maze_data[2999:2900] = maze_paths[29];
	assign maze_data[3099:3000]   = maze_paths[30];
	assign maze_data[3199:3100] = maze_paths[31];
	assign maze_data[3299:3200] = maze_paths[32];
	assign maze_data[3399:3300] = maze_paths[33];
	assign maze_data[3499:3400] = maze_paths[34];
	assign maze_data[3599:3500] = maze_paths[35];
	assign maze_data[3699:3600] = maze_paths[36];
	assign maze_data[3799:3700] = maze_paths[37];
	assign maze_data[3899:3800] = maze_paths[38];
	assign maze_data[3999:3900] = maze_paths[39];
	assign maze_data[4099:4000]   = maze_paths[40];
	assign maze_data[4199:4100] = maze_paths[41];
	assign maze_data[4299:4200] = maze_paths[42];
	assign maze_data[4399:4300] = maze_paths[43];
	assign maze_data[4499:4400] = maze_paths[44];
	assign maze_data[4599:4500] = maze_paths[45];
	assign maze_data[4699:4600] = maze_paths[46];
	assign maze_data[4799:4700] = maze_paths[47];
	assign maze_data[4899:4800] = maze_paths[48];
	assign maze_data[4999:4900] = maze_paths[49];
	assign maze_data[5099:5000]   = maze_paths[50];
	assign maze_data[5199:5100] = maze_paths[51];
	assign maze_data[5299:5200] = maze_paths[52];
	assign maze_data[5399:5300] = maze_paths[53];
	assign maze_data[5499:5400] = maze_paths[54];
	assign maze_data[5599:5500] = maze_paths[55];
	assign maze_data[5699:5600] = maze_paths[56];
	assign maze_data[5799:5700] = maze_paths[57];
	assign maze_data[5899:5800] = maze_paths[58];
	assign maze_data[5999:5900] = maze_paths[59];
	assign maze_data[6099:6000]   = maze_paths[60];
	assign maze_data[6199:6100] = maze_paths[61];
	assign maze_data[6299:6200] = maze_paths[62];
	assign maze_data[6399:6300] = maze_paths[63];
	assign maze_data[6499:6400] = maze_paths[64];
	assign maze_data[6599:6500] = maze_paths[65];
	assign maze_data[6699:6600] = maze_paths[66];
	assign maze_data[6799:6700] = maze_paths[67];
	assign maze_data[6899:6800] = maze_paths[68];
	assign maze_data[6999:6900] = maze_paths[69];
	assign maze_data[7099:7000]   = maze_paths[70];
	assign maze_data[7199:7100] = maze_paths[71];
	assign maze_data[7299:7200] = maze_paths[72];
	assign maze_data[7399:7300] = maze_paths[73];
	assign maze_data[7499:7400] = maze_paths[74];
	assign maze_data[7599:7500] = maze_paths[75];
	assign maze_data[7699:7600] = maze_paths[76];
	assign maze_data[7799:7700] = maze_paths[77];
	assign maze_data[7899:7800] = maze_paths[78];
	assign maze_data[7999:7900] = maze_paths[79];
	assign maze_data[8099:8000]   = maze_paths[80];
	assign maze_data[8199:8100] = maze_paths[81];
	assign maze_data[8299:8200] = maze_paths[82];
	assign maze_data[8399:8300] = maze_paths[83];
	assign maze_data[8499:8400] = maze_paths[84];
	assign maze_data[8599:8500] = maze_paths[85];
	assign maze_data[8699:8600] = maze_paths[86];
	assign maze_data[8799:8700] = maze_paths[87];
	assign maze_data[8899:8800] = maze_paths[88];
	assign maze_data[8999:8900] = maze_paths[89];
	assign maze_data[9099:9000]   = maze_paths[90];
	assign maze_data[9199:9100] = maze_paths[91];
	assign maze_data[9299:9200] = maze_paths[92];
	assign maze_data[9399:9300] = maze_paths[93];
	assign maze_data[9499:9400] = maze_paths[94];
	assign maze_data[9599:9500] = maze_paths[95];
	assign maze_data[9699:9600] = maze_paths[96];
	assign maze_data[9799:9700] = maze_paths[97];
	assign maze_data[9899:9800] = maze_paths[98];
	assign maze_data[9999:9900] = maze_paths[99];

endmodule
*/
/*	initial begin
		maze_paths [0] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [1] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [2] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [3] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [4] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [5] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [6] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [7] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [8] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [9] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [10] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [11] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [12] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [13] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [14] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [15] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [16] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [17] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [18] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [19] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [20] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [21] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [22] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [23] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [24] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [25] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [26] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [27] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [28] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [29] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [30] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [31] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [32] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [33] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [34] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [35] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [36] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [37] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [38] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [39] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [40] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [41] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [42] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [43] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [44] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [45] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [46] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [47] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [48] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [49] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [50] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [51] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [52] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [53] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [54] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [55] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [56] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [57] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [58] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [59] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [60] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [61] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [62] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [63] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [64] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [65] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [66] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [67] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [68] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [69] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [70] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [71] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [72] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [73] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [74] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [75] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [76] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [77] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [78] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [79] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [80] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [81] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [82] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [83] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [84] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [85] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [86] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [87] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [88] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [89] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [90] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [91] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [92] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [93] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [94] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
		maze_paths [95] <= 100'b0111010010011101001001110100100111010010011101001001110100100111010010011101001001110100100111010010;
		maze_paths [96] <= 100'b0000011111000001111100000111110000011111000001111100000111110000011111000001111100000111110000011111;
		maze_paths [97] <= 100'b0101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
		maze_paths [98] <= 100'b1100011011110001101111000110111100011011110001101111000110111100011011110001101111000110111100011011;
		maze_paths [99] <= 100'b1010101000101010100010101010001010101000101010100010101010001010101000101010100010101010001010101000;
*/