
module maze_carver
	(
		input clk,
		input start,
		input wire [2:0] x_dimension,
		input wire [2:0] y_dimension,
		output reg [64*64-1:0] maze_data,
		output reg finish
	);
	
	reg [15:0] i;
	reg [15:0] j;

	initial begin
		for (i = 0; i < 64; i = i + 1)
			for (j = 0; j < 64; j = j + 1)
				maze_data [i + 64*j] = 1;
//		maze_data = 4096'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
//		maze_data = 4096'b1011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010101101101001011010110110100101011011010010110101101101001011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110101010010110011010101010101000000101011011010101001011001101010101010100000010101101101010100101100110101010101010000001010110110101010010110011010101010101000001101010101010100000010101101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101101101001011010110110100101101011011010010110101011011011010110110101010010110011010101010101000001101010101010100000010101101101010100010101010111010101001011001101010101010100000110110101010010110011010101010101000001101101010100101100110101010101010000011011010101001011001101010101010100000110010011010100110011010010101101001010101011010100101011011011010110110101010010110011010101010101000001101010101010100000010101101101010100010101010101001101010011001101001010110100101010101101010010110110100101101011011010101001011001101010101010100000010101101101010100101100110101010101010000001010110110101010010110011010101010101000000010100000110101010101010000001010110110110101101101010100101100110101010101010000011010101010101000000101011011010101000101010101010011010100110011010010101101001010101011010100110011010010101101001010101011010100110111;
		maze_data = 4096'b1010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101101010101110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010110101010111010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101011010101010101010010101010101010110101010101010100101010101010101101010101010101001010101010101011;
		
	end
	
endmodule
